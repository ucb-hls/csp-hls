// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 5.1 (http://legupcomputing.com)
// Copyright (c) 2015-2017 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Tue Dec 12 00:21:01 2017
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This is a relative path to the directories where simulation and FPGA vendors' synthesis flow will run.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val,
	auto_pthread_wrapper_start,
	auto_pthread_wrapper_threadID,
	auto_pthread_wrapper_OC_1_start,
	auto_pthread_wrapper_OC_1_threadID,
	main_0_1_ready_from_sink,
	main_0_1_valid_to_sink,
	main_0_1_data_to_sink,
	main_0_3_ready_to_source,
	main_0_3_valid_from_source,
	main_0_3_data_from_source
);

parameter [4:0] LEGUP_0 = 5'd0;
parameter [4:0] LEGUP_F_main_BB__0_1 = 5'd1;
parameter [4:0] LEGUP_F_main_BB__0_2 = 5'd2;
parameter [4:0] LEGUP_F_main_BB__0_3 = 5'd3;
parameter [4:0] LEGUP_F_main_BB__0_4 = 5'd4;
parameter [4:0] LEGUP_F_main_BB__0_5 = 5'd5;
parameter [4:0] LEGUP_F_main_BB__0_6 = 5'd6;
parameter [4:0] LEGUP_F_main_BB__0_7 = 5'd7;
parameter [4:0] LEGUP_F_main_BB__0_8 = 5'd8;
parameter [4:0] LEGUP_F_main_BB__0_9 = 5'd9;
parameter [4:0] LEGUP_F_main_BB__0_10 = 5'd10;
parameter [4:0] LEGUP_F_main_BB__0_12 = 5'd12;
parameter [4:0] LEGUP_F_main_BB__0_14 = 5'd14;
parameter [4:0] LEGUP_F_main_BB__0_15 = 5'd15;
parameter [4:0] LEGUP_F_main_BB__0_16 = 5'd16;
parameter [4:0] LEGUP_F_main_BB__0_17 = 5'd17;
parameter [4:0] LEGUP_F_main_BB__0_18 = 5'd18;
parameter [4:0] LEGUP_F_main_BB__0_19 = 5'd19;
parameter [4:0] LEGUP_F_main_BB__0_20 = 5'd20;
parameter [4:0] LEGUP_F_main_BB__0_21 = 5'd21;
parameter [4:0] LEGUP_F_main_BB__0_22 = 5'd22;
parameter [4:0] LEGUP_F_main_BB__0_23 = 5'd23;
parameter [4:0] LEGUP_function_call_11 = 5'd11;
parameter [4:0] LEGUP_function_call_13 = 5'd13;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
output reg  auto_pthread_wrapper_start;
output reg [15:0] auto_pthread_wrapper_threadID;
output reg  auto_pthread_wrapper_OC_1_start;
output reg [15:0] auto_pthread_wrapper_OC_1_threadID;
input  main_0_1_ready_from_sink;
output reg  main_0_1_valid_to_sink;
output reg [63:0] main_0_1_data_to_sink;
output reg  main_0_3_ready_to_source;
input  main_0_3_valid_from_source;
input [63:0] main_0_3_data_from_source;
reg [4:0] cur_state;
reg [4:0] next_state;
reg  fsm_stall;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_enable_cond_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_not_accessed_due_to_stall_a;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_stalln_reg;
reg  main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_enable_cond_a;
reg  main_0_3_inputFIFO_consumed_valid;
reg  main_0_3_inputFIFO_consumed_taken;


always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  // synthesis parallel_case  
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB__0_1;
LEGUP_F_main_BB__0_1:
		next_state = LEGUP_F_main_BB__0_2;
LEGUP_F_main_BB__0_10:
		next_state = LEGUP_function_call_11;
LEGUP_F_main_BB__0_12:
		next_state = LEGUP_function_call_13;
LEGUP_F_main_BB__0_14:
		next_state = LEGUP_F_main_BB__0_15;
LEGUP_F_main_BB__0_15:
		next_state = LEGUP_F_main_BB__0_16;
LEGUP_F_main_BB__0_16:
		next_state = LEGUP_F_main_BB__0_17;
LEGUP_F_main_BB__0_17:
		next_state = LEGUP_F_main_BB__0_18;
LEGUP_F_main_BB__0_18:
		next_state = LEGUP_F_main_BB__0_19;
LEGUP_F_main_BB__0_19:
		next_state = LEGUP_F_main_BB__0_20;
LEGUP_F_main_BB__0_2:
		next_state = LEGUP_F_main_BB__0_3;
LEGUP_F_main_BB__0_20:
		next_state = LEGUP_F_main_BB__0_21;
LEGUP_F_main_BB__0_21:
		next_state = LEGUP_F_main_BB__0_22;
LEGUP_F_main_BB__0_22:
		next_state = LEGUP_F_main_BB__0_23;
LEGUP_F_main_BB__0_23:
		next_state = LEGUP_0;
LEGUP_F_main_BB__0_3:
		next_state = LEGUP_F_main_BB__0_4;
LEGUP_F_main_BB__0_4:
		next_state = LEGUP_F_main_BB__0_5;
LEGUP_F_main_BB__0_5:
		next_state = LEGUP_F_main_BB__0_6;
LEGUP_F_main_BB__0_6:
		next_state = LEGUP_F_main_BB__0_7;
LEGUP_F_main_BB__0_7:
		next_state = LEGUP_F_main_BB__0_8;
LEGUP_F_main_BB__0_8:
		next_state = LEGUP_F_main_BB__0_9;
LEGUP_F_main_BB__0_9:
		next_state = LEGUP_F_main_BB__0_10;
LEGUP_function_call_11:
		next_state = LEGUP_F_main_BB__0_12;
LEGUP_function_call_13:
		next_state = LEGUP_F_main_BB__0_14;
default:
	next_state = cur_state;
endcase

end
always @(*) begin
	fsm_stall = 1'd0;
	if (((cur_state == LEGUP_F_main_BB__0_1) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_2) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_3) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_4) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_5) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_6) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_7) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_8) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_9) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_10) & ~(main_0_1_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_14) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_15) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_16) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_17) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_18) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_19) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_20) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_21) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_22) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_main_BB__0_23) & ~(main_0_3_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_1) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_2) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_3) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_4) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_5) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_6) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_7) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_8) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_9) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_stalln_reg));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_1_valid_to_sink) & ~(main_0_1_ready_from_sink));
end
always @(posedge clk) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_enable_cond_a = ((cur_state == LEGUP_F_main_BB__0_10) & (main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_not_accessed_due_to_stall_a | main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_stalln_reg));
end
always @(posedge clk) begin
	if (main_0_3_inputFIFO_consumed_taken) begin
		main_0_3_inputFIFO_consumed_valid <= 1'd0;
	end
	if ((main_0_3_ready_to_source & main_0_3_valid_from_source)) begin
		main_0_3_inputFIFO_consumed_valid <= 1'd1;
	end
	if (reset) begin
		main_0_3_inputFIFO_consumed_valid <= 1'd0;
	end
end
always @(*) begin
	main_0_3_inputFIFO_consumed_taken = 1'd0;
	if (reset) begin
		main_0_3_inputFIFO_consumed_taken = 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB__0_14)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_15)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_16)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_17)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_18)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_19)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_20)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_21)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_22)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_main_BB__0_23)) begin
		main_0_3_inputFIFO_consumed_taken = ~(fsm_stall);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	/* main: %0*/
	/*   ret i32 0, !dbg !263, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_23)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	/* main: %0*/
	/*   ret i32 0, !dbg !263, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_23)) begin
		return_val <= 32'd0;
	end
end
always @(posedge clk) begin
	if (reset) begin
		auto_pthread_wrapper_start <= 1'd0;
	end
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper(%struct.FIFO* %1, %struct.FIFO* %2) #8, !dbg !235, !PTHREADNAME !237, !NUMTHREADS !238, !FUNCTIONID !202, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_10)) begin
		auto_pthread_wrapper_start <= 1'd1;
	end
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper(%struct.FIFO* %1, %struct.FIFO* %2) #8, !dbg !235, !PTHREADNAME !237, !NUMTHREADS !238, !FUNCTIONID !202, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if (((cur_state == LEGUP_function_call_11) & ~(fsm_stall))) begin
		auto_pthread_wrapper_start <= 1'd0;
	end
end
always @(posedge clk) begin
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper(%struct.FIFO* %1, %struct.FIFO* %2) #8, !dbg !235, !PTHREADNAME !237, !NUMTHREADS !238, !FUNCTIONID !202, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_10)) begin
		auto_pthread_wrapper_threadID <= 1'd0;
	end
end
always @(posedge clk) begin
	if (reset) begin
		auto_pthread_wrapper_OC_1_start <= 1'd0;
	end
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper_OC_1(%struct.FIFO* %2, %struct.FIFO* %3) #8, !dbg !240, !PTHREADNAME !241, !NUMTHREADS !238, !FUNCTIONID !238, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_12)) begin
		auto_pthread_wrapper_OC_1_start <= 1'd1;
	end
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper_OC_1(%struct.FIFO* %2, %struct.FIFO* %3) #8, !dbg !240, !PTHREADNAME !241, !NUMTHREADS !238, !FUNCTIONID !238, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if (((cur_state == LEGUP_function_call_13) & ~(fsm_stall))) begin
		auto_pthread_wrapper_OC_1_start <= 1'd0;
	end
end
always @(posedge clk) begin
	/* main: %0*/
	/*   call fastcc void @auto_pthread_wrapper_OC_1(%struct.FIFO* %2, %struct.FIFO* %3) #8, !dbg !240, !PTHREADNAME !241, !NUMTHREADS !238, !FUNCTIONID !238, !TYPE !239, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_12)) begin
		auto_pthread_wrapper_OC_1_threadID <= 1'd0;
	end
end
always @(*) begin
	main_0_1_valid_to_sink = 1'd0;
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_1_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_2_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_3_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_4_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_5_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_6_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_7_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_8_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_9_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
	if (main_0_1_outputFIFO_LEGUP_F_main_BB__0_10_enable_cond_a) begin
		main_0_1_valid_to_sink = 1'd1;
	end
end
always @(*) begin
	main_0_1_data_to_sink = 64'd0;
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 0) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_1)) begin
		main_0_1_data_to_sink = 64'd0;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 1) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_2)) begin
		main_0_1_data_to_sink = 64'd1;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 4) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_3)) begin
		main_0_1_data_to_sink = 64'd4;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 9) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_4)) begin
		main_0_1_data_to_sink = 64'd9;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 16) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_5)) begin
		main_0_1_data_to_sink = 64'd16;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 25) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_6)) begin
		main_0_1_data_to_sink = 64'd25;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 36) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_7)) begin
		main_0_1_data_to_sink = 64'd36;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 49) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_8)) begin
		main_0_1_data_to_sink = 64'd49;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 64) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_9)) begin
		main_0_1_data_to_sink = 64'd64;
	end
	/* main: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %1, i64 81) #7, !dbg !226, !MSB !201, !LSB !202, !extendFrom !201*/
	if ((cur_state == LEGUP_F_main_BB__0_10)) begin
		main_0_1_data_to_sink = 64'd81;
	end
end
always @(*) begin
	main_0_3_ready_to_source = (~(main_0_3_inputFIFO_consumed_valid) | main_0_3_inputFIFO_consumed_taken);
	if (reset) begin
		main_0_3_ready_to_source = 1'd0;
	end
end

endmodule
`timescale 1 ns / 1 ns
module auto_pthread_wrapper
(
	clk,
	reset,
	start,
	finish,
	main_0_1_ready_to_source,
	main_0_1_valid_from_source,
	main_0_1_data_from_source,
	main_0_2_ready_from_sink,
	main_0_2_valid_to_sink,
	main_0_2_data_to_sink
);

parameter [3:0] LEGUP_0 = 4'd0;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_1 = 4'd1;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_2 = 4'd2;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_3 = 4'd3;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_4 = 4'd4;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_5 = 4'd5;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_6 = 4'd6;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_7 = 4'd7;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_8 = 4'd8;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_9 = 4'd9;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_10 = 4'd10;
parameter [3:0] LEGUP_F_auto_pthread_wrapper_BB__0_11 = 4'd11;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg  main_0_1_ready_to_source;
input  main_0_1_valid_from_source;
input [63:0] main_0_1_data_from_source;
input  main_0_2_ready_from_sink;
output reg  main_0_2_valid_to_sink;
output reg [63:0] main_0_2_data_to_sink;
reg [3:0] cur_state;
reg [3:0] next_state;
reg  fsm_stall;
reg [62:0] auto_pthread_wrapper_0_1;
reg [63:0] auto_pthread_wrapper_0_2;
reg [63:0] auto_pthread_wrapper_0_3;
reg [63:0] auto_pthread_wrapper_0_3_reg;
reg [62:0] auto_pthread_wrapper_0_4;
reg [63:0] auto_pthread_wrapper_0_5;
reg [63:0] auto_pthread_wrapper_0_6;
reg [63:0] auto_pthread_wrapper_0_6_reg;
reg [62:0] auto_pthread_wrapper_0_7;
reg [63:0] auto_pthread_wrapper_0_8;
reg [63:0] auto_pthread_wrapper_0_9;
reg [63:0] auto_pthread_wrapper_0_9_reg;
reg [62:0] auto_pthread_wrapper_0_10;
reg [63:0] auto_pthread_wrapper_0_11;
reg [63:0] auto_pthread_wrapper_0_12;
reg [63:0] auto_pthread_wrapper_0_12_reg;
reg [62:0] auto_pthread_wrapper_0_13;
reg [63:0] auto_pthread_wrapper_0_14;
reg [63:0] auto_pthread_wrapper_0_15;
reg [63:0] auto_pthread_wrapper_0_15_reg;
reg [62:0] auto_pthread_wrapper_0_16;
reg [63:0] auto_pthread_wrapper_0_17;
reg [63:0] auto_pthread_wrapper_0_18;
reg [63:0] auto_pthread_wrapper_0_18_reg;
reg [62:0] auto_pthread_wrapper_0_19;
reg [63:0] auto_pthread_wrapper_0_20;
reg [63:0] auto_pthread_wrapper_0_21;
reg [63:0] auto_pthread_wrapper_0_21_reg;
reg [62:0] auto_pthread_wrapper_0_22;
reg [63:0] auto_pthread_wrapper_0_23;
reg [63:0] auto_pthread_wrapper_0_24;
reg [63:0] auto_pthread_wrapper_0_24_reg;
reg [62:0] auto_pthread_wrapper_0_25;
reg [63:0] auto_pthread_wrapper_0_26;
reg [63:0] auto_pthread_wrapper_0_27;
reg [63:0] auto_pthread_wrapper_0_27_reg;
reg [62:0] auto_pthread_wrapper_0_28;
reg [63:0] auto_pthread_wrapper_0_29;
reg [63:0] auto_pthread_wrapper_0_30;
reg [63:0] auto_pthread_wrapper_0_30_reg;
reg  main_0_1_inputFIFO_consumed_valid;
reg [63:0] main_0_1_inputFIFO_consumed_data;
reg  main_0_1_inputFIFO_consumed_taken;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_enable_cond_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_not_accessed_due_to_stall_a;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_stalln_reg;
reg  main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_enable_cond_a;


always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  // synthesis parallel_case  
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_1;
LEGUP_F_auto_pthread_wrapper_BB__0_1:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_2;
LEGUP_F_auto_pthread_wrapper_BB__0_10:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_11;
LEGUP_F_auto_pthread_wrapper_BB__0_11:
		next_state = LEGUP_0;
LEGUP_F_auto_pthread_wrapper_BB__0_2:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_3;
LEGUP_F_auto_pthread_wrapper_BB__0_3:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_4;
LEGUP_F_auto_pthread_wrapper_BB__0_4:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_5;
LEGUP_F_auto_pthread_wrapper_BB__0_5:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_6;
LEGUP_F_auto_pthread_wrapper_BB__0_6:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_7;
LEGUP_F_auto_pthread_wrapper_BB__0_7:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_8;
LEGUP_F_auto_pthread_wrapper_BB__0_8:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_9;
LEGUP_F_auto_pthread_wrapper_BB__0_9:
		next_state = LEGUP_F_auto_pthread_wrapper_BB__0_10;
default:
	next_state = cur_state;
endcase

end
always @(*) begin
	fsm_stall = 1'd0;
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_1) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10) & ~(main_0_1_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_11) & ~(main_0_2_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_1 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %2 = shl i64 %1, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_2 = ({1'd0,auto_pthread_wrapper_0_1} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %3 = or i64 %2, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_3 = (auto_pthread_wrapper_0_2 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %3 = or i64 %2, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_1)) begin
		auto_pthread_wrapper_0_3_reg <= auto_pthread_wrapper_0_3;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_4 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %5 = shl i64 %4, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_5 = ({1'd0,auto_pthread_wrapper_0_4} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %6 = or i64 %5, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_6 = (auto_pthread_wrapper_0_5 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %6 = or i64 %5, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2)) begin
		auto_pthread_wrapper_0_6_reg <= auto_pthread_wrapper_0_6;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_7 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %8 = shl i64 %7, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_8 = ({1'd0,auto_pthread_wrapper_0_7} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %9 = or i64 %8, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_9 = (auto_pthread_wrapper_0_8 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %9 = or i64 %8, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3)) begin
		auto_pthread_wrapper_0_9_reg <= auto_pthread_wrapper_0_9;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_10 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %11 = shl i64 %10, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_11 = ({1'd0,auto_pthread_wrapper_0_10} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %12 = or i64 %11, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_12 = (auto_pthread_wrapper_0_11 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %12 = or i64 %11, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4)) begin
		auto_pthread_wrapper_0_12_reg <= auto_pthread_wrapper_0_12;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_13 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %14 = shl i64 %13, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_14 = ({1'd0,auto_pthread_wrapper_0_13} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %15 = or i64 %14, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_15 = (auto_pthread_wrapper_0_14 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %15 = or i64 %14, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5)) begin
		auto_pthread_wrapper_0_15_reg <= auto_pthread_wrapper_0_15;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_16 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %17 = shl i64 %16, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_17 = ({1'd0,auto_pthread_wrapper_0_16} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %18 = or i64 %17, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_18 = (auto_pthread_wrapper_0_17 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %18 = or i64 %17, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6)) begin
		auto_pthread_wrapper_0_18_reg <= auto_pthread_wrapper_0_18;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_19 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %20 = shl i64 %19, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_20 = ({1'd0,auto_pthread_wrapper_0_19} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %21 = or i64 %20, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_21 = (auto_pthread_wrapper_0_20 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %21 = or i64 %20, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7)) begin
		auto_pthread_wrapper_0_21_reg <= auto_pthread_wrapper_0_21;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_22 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %23 = shl i64 %22, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_23 = ({1'd0,auto_pthread_wrapper_0_22} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %24 = or i64 %23, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_24 = (auto_pthread_wrapper_0_23 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %24 = or i64 %23, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8)) begin
		auto_pthread_wrapper_0_24_reg <= auto_pthread_wrapper_0_24;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_25 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %26 = shl i64 %25, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_26 = ({1'd0,auto_pthread_wrapper_0_25} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %27 = or i64 %26, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_27 = (auto_pthread_wrapper_0_26 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %27 = or i64 %26, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9)) begin
		auto_pthread_wrapper_0_27_reg <= auto_pthread_wrapper_0_27;
	end
end
always @(*) begin
	auto_pthread_wrapper_0_28 = main_0_1_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %29 = shl i64 %28, 1, !dbg !302, !MSB !303, !LSB !304, !extendFrom !303*/
		auto_pthread_wrapper_0_29 = ({1'd0,auto_pthread_wrapper_0_28} <<< (64'd1 % 64'd64));
end
always @(*) begin
	/* auto_pthread_wrapper: %0*/
	/*   %30 = or i64 %29, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
		auto_pthread_wrapper_0_30 = (auto_pthread_wrapper_0_29 | 64'd1);
end
always @(posedge clk) begin
	/* auto_pthread_wrapper: %0*/
	/*   %30 = or i64 %29, 1, !dbg !316, !MSB !303, !LSB !256, !extendFrom !303*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10)) begin
		auto_pthread_wrapper_0_30_reg <= auto_pthread_wrapper_0_30;
	end
end
always @(posedge clk) begin
	if (main_0_1_inputFIFO_consumed_taken) begin
		main_0_1_inputFIFO_consumed_valid <= 1'd0;
	end
	if ((main_0_1_ready_to_source & main_0_1_valid_from_source)) begin
		main_0_1_inputFIFO_consumed_valid <= 1'd1;
	end
	if (reset) begin
		main_0_1_inputFIFO_consumed_valid <= 1'd0;
	end
end
always @(posedge clk) begin
	if ((main_0_1_ready_to_source & main_0_1_valid_from_source)) begin
		main_0_1_inputFIFO_consumed_data <= main_0_1_data_from_source;
	end
	if (reset) begin
		main_0_1_inputFIFO_consumed_data <= 1'd0;
	end
end
always @(*) begin
	main_0_1_inputFIFO_consumed_taken = 1'd0;
	if (reset) begin
		main_0_1_inputFIFO_consumed_taken = 1'd0;
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_1)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10)) begin
		main_0_1_inputFIFO_consumed_taken = ~(fsm_stall);
	end
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_stalln_reg));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_2_valid_to_sink) & ~(main_0_2_ready_from_sink));
end
always @(posedge clk) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_11) & (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_not_accessed_due_to_stall_a | main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_stalln_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	/* auto_pthread_wrapper: %0*/
	/*   ret void, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_11)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(*) begin
	main_0_1_ready_to_source = (~(main_0_1_inputFIFO_consumed_valid) | main_0_1_inputFIFO_consumed_taken);
	if (reset) begin
		main_0_1_ready_to_source = 1'd0;
	end
end
always @(*) begin
	main_0_2_valid_to_sink = 1'd0;
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_2_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_3_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_4_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_5_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_6_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_7_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_8_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_9_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_10_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
	if (main_0_2_outputFIFO_LEGUP_F_auto_pthread_wrapper_BB__0_11_enable_cond_a) begin
		main_0_2_valid_to_sink = 1'd1;
	end
end
always @(*) begin
	main_0_2_data_to_sink = 64'd0;
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %3) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_2)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_3_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %6) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_3)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_6_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %9) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_4)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_9_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %12) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_5)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_12_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %15) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_6)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_15_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %18) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_7)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_18_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %21) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_8)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_21_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %24) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_9)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_24_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %27) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_10)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_27_reg;
	end
	/* auto_pthread_wrapper: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %30) #7, !dbg !319, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_BB__0_11)) begin
		main_0_2_data_to_sink = auto_pthread_wrapper_0_30_reg;
	end
end

endmodule
`timescale 1 ns / 1 ns
module auto_pthread_wrapper_OC_1
(
	clk,
	reset,
	start,
	finish,
	main_0_2_ready_to_source,
	main_0_2_valid_from_source,
	main_0_2_data_from_source,
	main_0_3_ready_from_sink,
	main_0_3_valid_to_sink,
	main_0_3_data_to_sink
);

parameter [6:0] LEGUP_0 = 7'd0;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1 = 7'd1;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2 = 7'd2;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3 = 7'd3;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4 = 7'd4;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5 = 7'd5;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6 = 7'd6;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7 = 7'd7;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8 = 7'd8;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9 = 7'd9;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10 = 7'd10;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_11 = 7'd11;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_12 = 7'd12;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_13 = 7'd13;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_14 = 7'd14;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_15 = 7'd15;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_16 = 7'd16;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_17 = 7'd17;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_18 = 7'd18;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_19 = 7'd19;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_20 = 7'd20;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_21 = 7'd21;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_22 = 7'd22;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_23 = 7'd23;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_24 = 7'd24;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_25 = 7'd25;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_26 = 7'd26;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_27 = 7'd27;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_28 = 7'd28;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_29 = 7'd29;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_30 = 7'd30;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_31 = 7'd31;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_32 = 7'd32;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_33 = 7'd33;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_34 = 7'd34;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_35 = 7'd35;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_36 = 7'd36;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_37 = 7'd37;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_38 = 7'd38;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_39 = 7'd39;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_40 = 7'd40;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_41 = 7'd41;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_42 = 7'd42;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_43 = 7'd43;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_44 = 7'd44;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_45 = 7'd45;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_46 = 7'd46;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_47 = 7'd47;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_48 = 7'd48;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_49 = 7'd49;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_50 = 7'd50;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_51 = 7'd51;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_52 = 7'd52;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_53 = 7'd53;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_54 = 7'd54;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_55 = 7'd55;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_56 = 7'd56;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_57 = 7'd57;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_58 = 7'd58;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_59 = 7'd59;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_60 = 7'd60;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_61 = 7'd61;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_62 = 7'd62;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_63 = 7'd63;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_64 = 7'd64;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65 = 7'd65;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66 = 7'd66;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67 = 7'd67;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68 = 7'd68;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69 = 7'd69;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70 = 7'd70;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71 = 7'd71;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72 = 7'd72;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73 = 7'd73;
parameter [6:0] LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74 = 7'd74;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg  main_0_2_ready_to_source;
input  main_0_2_valid_from_source;
input [63:0] main_0_2_data_from_source;
input  main_0_3_ready_from_sink;
output reg  main_0_3_valid_to_sink;
output reg [63:0] main_0_3_data_to_sink;
reg [6:0] cur_state;
reg [6:0] next_state;
reg  fsm_stall;
reg [63:0] auto_pthread_wrapper_OC_1_0_1;
reg [63:0] auto_pthread_wrapper_OC_1_0_2;
reg [62:0] auto_pthread_wrapper_OC_1_0_3;
reg [63:0] auto_pthread_wrapper_OC_1_0_4;
reg [63:0] auto_pthread_wrapper_OC_1_0_5;
reg [62:0] auto_pthread_wrapper_OC_1_0_6;
reg [63:0] auto_pthread_wrapper_OC_1_0_7;
reg [63:0] auto_pthread_wrapper_OC_1_0_8;
reg [62:0] auto_pthread_wrapper_OC_1_0_9;
reg [63:0] auto_pthread_wrapper_OC_1_0_10;
reg [63:0] auto_pthread_wrapper_OC_1_0_11;
reg [62:0] auto_pthread_wrapper_OC_1_0_12;
reg [63:0] auto_pthread_wrapper_OC_1_0_13;
reg [63:0] auto_pthread_wrapper_OC_1_0_14;
reg [62:0] auto_pthread_wrapper_OC_1_0_15;
reg [63:0] auto_pthread_wrapper_OC_1_0_16;
reg [63:0] auto_pthread_wrapper_OC_1_0_17;
reg [62:0] auto_pthread_wrapper_OC_1_0_18;
reg [63:0] auto_pthread_wrapper_OC_1_0_19;
reg [63:0] auto_pthread_wrapper_OC_1_0_20;
reg [62:0] auto_pthread_wrapper_OC_1_0_21;
reg [63:0] auto_pthread_wrapper_OC_1_0_22;
reg [63:0] auto_pthread_wrapper_OC_1_0_23;
reg [62:0] auto_pthread_wrapper_OC_1_0_24;
reg [63:0] auto_pthread_wrapper_OC_1_0_25;
reg [63:0] auto_pthread_wrapper_OC_1_0_26;
reg [62:0] auto_pthread_wrapper_OC_1_0_27;
reg [63:0] auto_pthread_wrapper_OC_1_0_28;
reg [63:0] auto_pthread_wrapper_OC_1_0_29;
reg [62:0] auto_pthread_wrapper_OC_1_0_30;
reg [63:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_op0;
reg [3:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_op1;
reg  auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clock;
reg  auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_aclr;
reg  auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clken;
reg [63:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_numer;
reg [3:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_denom;
wire [63:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_quotient;
wire [3:0] auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_remain;
reg [63:0] divide_auto_pthread_wrapper_OC_1_0_3_temp_out;
reg  divide_auto_pthread_wrapper_OC_1_0_3_en;
reg [62:0] divide_auto_pthread_wrapper_OC_1_0_3_out;
reg [62:0] auto_pthread_wrapper_OC_1_signed_divide_64_0;
reg  main_0_2_inputFIFO_consumed_valid;
reg [63:0] main_0_2_inputFIFO_consumed_data;
reg  main_0_2_inputFIFO_consumed_taken;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_enable_cond_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_not_accessed_due_to_stall_a;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_stalln_reg;
reg  main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_enable_cond_a;

/*   %3 = sdiv i64 %2, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
lpm_divide auto_pthread_wrapper_OC_1_signed_divide_64_0_inst (
	.clock (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clock),
	.aclr (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_aclr),
	.clken (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clken),
	.numer (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_numer),
	.denom (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_denom),
	.quotient (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_quotient),
	.remain (auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_remain)
);

defparam
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_widthn = 64,
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_widthd = 4,
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_drepresentation = "SIGNED",
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_nrepresentation = "SIGNED",
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_hint = "LPM_REMAINDERPOSITIVE=FALSE",
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst.lpm_pipeline = 64;


always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  // synthesis parallel_case  
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_11;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_11:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_12;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_12:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_13;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_13:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_14;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_14:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_15;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_15:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_16;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_16:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_17;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_17:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_18;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_18:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_19;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_19:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_20;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_20:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_21;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_21:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_22;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_22:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_23;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_23:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_24;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_24:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_25;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_25:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_26;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_26:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_27;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_27:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_28;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_28:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_29;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_29:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_30;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_30:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_31;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_31:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_32;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_32:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_33;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_33:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_34;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_34:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_35;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_35:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_36;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_36:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_37;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_37:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_38;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_38:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_39;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_39:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_40;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_40:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_41;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_41:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_42;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_42:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_43;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_43:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_44;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_44:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_45;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_45:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_46;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_46:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_47;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_47:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_48;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_48:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_49;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_49:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_50;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_50:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_51;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_51:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_52;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_52:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_53;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_53:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_54;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_54:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_55;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_55:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_56;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_56:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_57;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_57:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_58;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_58:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_59;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_59:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_60;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_60:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_61;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_61:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_62;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_62:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_63;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_63:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_64;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_64:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74:
		next_state = LEGUP_0;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9;
LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9:
		next_state = LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10;
default:
	next_state = cur_state;
endcase

end
always @(*) begin
	fsm_stall = 1'd0;
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10) & ~(main_0_2_inputFIFO_consumed_valid))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
	if (((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74) & ~(main_0_3_ready_from_sink))) begin
		fsm_stall = 1'd1;
	end
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_1 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %2 = add i64 %1, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_2 = (auto_pthread_wrapper_OC_1_0_1 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_3 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_4 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %5 = add i64 %4, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_5 = (auto_pthread_wrapper_OC_1_0_4 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_6 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_7 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %8 = add i64 %7, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_8 = (auto_pthread_wrapper_OC_1_0_7 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_9 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_10 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %11 = add i64 %10, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_11 = (auto_pthread_wrapper_OC_1_0_10 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_12 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_13 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %14 = add i64 %13, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_14 = (auto_pthread_wrapper_OC_1_0_13 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_15 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_16 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %17 = add i64 %16, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_17 = (auto_pthread_wrapper_OC_1_0_16 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_18 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_19 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %20 = add i64 %19, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_20 = (auto_pthread_wrapper_OC_1_0_19 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_21 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_22 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %23 = add i64 %22, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_23 = (auto_pthread_wrapper_OC_1_0_22 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_24 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_25 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %26 = add i64 %25, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_26 = (auto_pthread_wrapper_OC_1_0_25 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_27 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_28 = main_0_2_inputFIFO_consumed_data;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %29 = add i64 %28, -1, !dbg !300, !MSB !284, !LSB !256, !extendFrom !284*/
		auto_pthread_wrapper_OC_1_0_29 = (auto_pthread_wrapper_OC_1_0_28 + $signed(-64'd1));
end
always @(*) begin
	auto_pthread_wrapper_OC_1_0_30 = auto_pthread_wrapper_OC_1_signed_divide_64_0;
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %3 = sdiv i64 %2, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %6 = sdiv i64 %5, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_5;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %9 = sdiv i64 %8, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_8;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %12 = sdiv i64 %11, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_11;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %15 = sdiv i64 %14, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_14;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %18 = sdiv i64 %17, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_17;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %21 = sdiv i64 %20, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_20;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %24 = sdiv i64 %23, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_23;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %27 = sdiv i64 %26, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_26;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %30 = sdiv i64 %29, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else /* if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10)) */ begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op0 = auto_pthread_wrapper_OC_1_0_29;
	end
end
always @(*) begin
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %3 = sdiv i64 %2, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %6 = sdiv i64 %5, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %9 = sdiv i64 %8, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %12 = sdiv i64 %11, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %15 = sdiv i64 %14, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %18 = sdiv i64 %17, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %21 = sdiv i64 %20, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %24 = sdiv i64 %23, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %27 = sdiv i64 %26, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9)) begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   %30 = sdiv i64 %29, 2, !dbg !312, !MSB !284, !LSB !256, !extendFrom !313*/
	else /* if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10)) */ begin
		auto_pthread_wrapper_OC_1_signed_divide_64_0_op1 = 64'd2;
	end
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clock = clk;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_aclr = reset;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_clken = divide_auto_pthread_wrapper_OC_1_0_3_en;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_numer = auto_pthread_wrapper_OC_1_signed_divide_64_0_op0;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_denom = auto_pthread_wrapper_OC_1_signed_divide_64_0_op1;
end
always @(*) begin
	divide_auto_pthread_wrapper_OC_1_0_3_temp_out = auto_pthread_wrapper_OC_1_signed_divide_64_0_inst_quotient;
end
always @(*) begin
	divide_auto_pthread_wrapper_OC_1_0_3_en = ~(fsm_stall);
end
always @(*) begin
	divide_auto_pthread_wrapper_OC_1_0_3_out = divide_auto_pthread_wrapper_OC_1_0_3_temp_out;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_signed_divide_64_0 = divide_auto_pthread_wrapper_OC_1_0_3_out;
end
always @(posedge clk) begin
	if (main_0_2_inputFIFO_consumed_taken) begin
		main_0_2_inputFIFO_consumed_valid <= 1'd0;
	end
	if ((main_0_2_ready_to_source & main_0_2_valid_from_source)) begin
		main_0_2_inputFIFO_consumed_valid <= 1'd1;
	end
	if (reset) begin
		main_0_2_inputFIFO_consumed_valid <= 1'd0;
	end
end
always @(posedge clk) begin
	if ((main_0_2_ready_to_source & main_0_2_valid_from_source)) begin
		main_0_2_inputFIFO_consumed_data <= main_0_2_data_from_source;
	end
	if (reset) begin
		main_0_2_inputFIFO_consumed_data <= 1'd0;
	end
end
always @(*) begin
	main_0_2_inputFIFO_consumed_taken = 1'd0;
	if (reset) begin
		main_0_2_inputFIFO_consumed_taken = 1'd0;
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_1)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_2)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_3)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_4)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_5)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_6)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_7)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_8)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_9)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_10)) begin
		main_0_2_inputFIFO_consumed_taken = ~(fsm_stall);
	end
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_stalln_reg));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_not_accessed_due_to_stall_a <= ((fsm_stall & main_0_3_valid_to_sink) & ~(main_0_3_ready_from_sink));
end
always @(posedge clk) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_stalln_reg <= ~(fsm_stall);
end
always @(*) begin
	main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_enable_cond_a = ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74) & (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_not_accessed_due_to_stall_a | main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_stalln_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   ret void, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(*) begin
	main_0_2_ready_to_source = (~(main_0_2_inputFIFO_consumed_valid) | main_0_2_inputFIFO_consumed_taken);
	if (reset) begin
		main_0_2_ready_to_source = 1'd0;
	end
end
always @(*) begin
	main_0_3_valid_to_sink = 1'd0;
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
	if (main_0_3_outputFIFO_LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74_enable_cond_a) begin
		main_0_3_valid_to_sink = 1'd1;
	end
end
always @(*) begin
	main_0_3_data_to_sink = 64'd0;
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %3) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_65)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_3[62]}},auto_pthread_wrapper_OC_1_0_3};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %6) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_66)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_6[62]}},auto_pthread_wrapper_OC_1_0_6};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %9) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_67)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_9[62]}},auto_pthread_wrapper_OC_1_0_9};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %12) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_68)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_12[62]}},auto_pthread_wrapper_OC_1_0_12};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %15) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_69)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_15[62]}},auto_pthread_wrapper_OC_1_0_15};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %18) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_70)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_18[62]}},auto_pthread_wrapper_OC_1_0_18};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %21) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_71)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_21[62]}},auto_pthread_wrapper_OC_1_0_21};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %24) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_72)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_24[62]}},auto_pthread_wrapper_OC_1_0_24};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %27) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_73)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_27[62]}},auto_pthread_wrapper_OC_1_0_27};
	end
	/* auto_pthread_wrapper_OC_1: %0*/
	/*   tail call void @fifo_write(%struct.FIFO* %.0.1.val, i64 %30) #7, !dbg !316, !MSB !255, !LSB !256, !extendFrom !255*/
	if ((cur_state == LEGUP_F_auto_pthread_wrapper_OC_1_BB__0_74)) begin
		main_0_3_data_to_sink = {{1{auto_pthread_wrapper_OC_1_0_30[62]}},auto_pthread_wrapper_OC_1_0_30};
	end
end

endmodule
`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
wire  main_inst_auto_pthread_wrapper_start;
wire [15:0] main_inst_auto_pthread_wrapper_threadID;
wire  main_inst_auto_pthread_wrapper_OC_1_start;
wire [15:0] main_inst_auto_pthread_wrapper_OC_1_threadID;
reg  main_inst_main_0_1_ready_from_sink;
wire  main_inst_main_0_1_valid_to_sink;
wire [63:0] main_inst_main_0_1_data_to_sink;
wire  main_inst_main_0_3_ready_to_source;
reg  main_inst_main_0_3_valid_from_source;
reg [63:0] main_inst_main_0_3_data_from_source;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;
reg  main_0_1_inst_clk;
reg  main_0_1_inst_reset;
reg  main_0_1_inst_clken;
reg  main_0_1_inst_write_en;
reg [63:0] main_0_1_inst_write_data;
reg  main_0_1_inst_read_en;
wire [63:0] main_0_1_inst_read_data;
wire  main_0_1_inst_full;
wire  main_0_1_inst_almost_full;
wire  main_0_1_inst_empty;
wire  main_0_1_inst_almost_empty;
wire [4:0] main_0_1_inst_usedw;
reg  main_0_3_inst_clk;
reg  main_0_3_inst_reset;
reg  main_0_3_inst_clken;
reg  main_0_3_inst_write_en;
reg [63:0] main_0_3_inst_write_data;
reg  main_0_3_inst_read_en;
wire [63:0] main_0_3_inst_read_data;
wire  main_0_3_inst_full;
wire  main_0_3_inst_almost_full;
wire  main_0_3_inst_empty;
wire  main_0_3_inst_almost_empty;
wire [4:0] main_0_3_inst_usedw;
reg  auto_pthread_wrapper_inst_clk;
reg  auto_pthread_wrapper_inst_reset;
reg  auto_pthread_wrapper_inst_start;
wire  auto_pthread_wrapper_inst_finish;
wire  auto_pthread_wrapper_inst_main_0_1_ready_to_source;
reg  auto_pthread_wrapper_inst_main_0_1_valid_from_source;
reg [63:0] auto_pthread_wrapper_inst_main_0_1_data_from_source;
reg  auto_pthread_wrapper_inst_main_0_2_ready_from_sink;
wire  auto_pthread_wrapper_inst_main_0_2_valid_to_sink;
wire [63:0] auto_pthread_wrapper_inst_main_0_2_data_to_sink;
reg  auto_pthread_wrapper_inst_finish_reg;
reg  main_0_2_inst_clk;
reg  main_0_2_inst_reset;
reg  main_0_2_inst_clken;
reg  main_0_2_inst_write_en;
reg [63:0] main_0_2_inst_write_data;
reg  main_0_2_inst_read_en;
wire [63:0] main_0_2_inst_read_data;
wire  main_0_2_inst_full;
wire  main_0_2_inst_almost_full;
wire  main_0_2_inst_empty;
wire  main_0_2_inst_almost_empty;
wire [4:0] main_0_2_inst_usedw;
reg  auto_pthread_wrapper_OC_1_inst_clk;
reg  auto_pthread_wrapper_OC_1_inst_reset;
reg  auto_pthread_wrapper_OC_1_inst_start;
wire  auto_pthread_wrapper_OC_1_inst_finish;
wire  auto_pthread_wrapper_OC_1_inst_main_0_2_ready_to_source;
reg  auto_pthread_wrapper_OC_1_inst_main_0_2_valid_from_source;
reg [63:0] auto_pthread_wrapper_OC_1_inst_main_0_2_data_from_source;
reg  auto_pthread_wrapper_OC_1_inst_main_0_3_ready_from_sink;
wire  auto_pthread_wrapper_OC_1_inst_main_0_3_valid_to_sink;
wire [63:0] auto_pthread_wrapper_OC_1_inst_main_0_3_data_to_sink;
reg  auto_pthread_wrapper_OC_1_inst_finish_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val),
	.auto_pthread_wrapper_start (main_inst_auto_pthread_wrapper_start),
	.auto_pthread_wrapper_threadID (main_inst_auto_pthread_wrapper_threadID),
	.auto_pthread_wrapper_OC_1_start (main_inst_auto_pthread_wrapper_OC_1_start),
	.auto_pthread_wrapper_OC_1_threadID (main_inst_auto_pthread_wrapper_OC_1_threadID),
	.main_0_1_ready_from_sink (main_inst_main_0_1_ready_from_sink),
	.main_0_1_valid_to_sink (main_inst_main_0_1_valid_to_sink),
	.main_0_1_data_to_sink (main_inst_main_0_1_data_to_sink),
	.main_0_3_ready_to_source (main_inst_main_0_3_ready_to_source),
	.main_0_3_valid_from_source (main_inst_main_0_3_valid_from_source),
	.main_0_3_data_from_source (main_inst_main_0_3_data_from_source)
);



fwft_fifo main_0_1_inst (
	.clk (main_0_1_inst_clk),
	.reset (main_0_1_inst_reset),
	.clken (main_0_1_inst_clken),
	.write_en (main_0_1_inst_write_en),
	.write_data (main_0_1_inst_write_data),
	.read_en (main_0_1_inst_read_en),
	.read_data (main_0_1_inst_read_data),
	.full (main_0_1_inst_full),
	.almost_full (main_0_1_inst_almost_full),
	.empty (main_0_1_inst_empty),
	.almost_empty (main_0_1_inst_almost_empty),
	.usedw (main_0_1_inst_usedw)
);

defparam
	main_0_1_inst.width = 64,
	main_0_1_inst.depth = 10,
	main_0_1_inst.widthad = 4;


fwft_fifo main_0_3_inst (
	.clk (main_0_3_inst_clk),
	.reset (main_0_3_inst_reset),
	.clken (main_0_3_inst_clken),
	.write_en (main_0_3_inst_write_en),
	.write_data (main_0_3_inst_write_data),
	.read_en (main_0_3_inst_read_en),
	.read_data (main_0_3_inst_read_data),
	.full (main_0_3_inst_full),
	.almost_full (main_0_3_inst_almost_full),
	.empty (main_0_3_inst_empty),
	.almost_empty (main_0_3_inst_almost_empty),
	.usedw (main_0_3_inst_usedw)
);

defparam
	main_0_3_inst.width = 64,
	main_0_3_inst.depth = 10,
	main_0_3_inst.widthad = 4;


auto_pthread_wrapper auto_pthread_wrapper_inst (
	.clk (auto_pthread_wrapper_inst_clk),
	.reset (auto_pthread_wrapper_inst_reset),
	.start (auto_pthread_wrapper_inst_start),
	.finish (auto_pthread_wrapper_inst_finish),
	.main_0_1_ready_to_source (auto_pthread_wrapper_inst_main_0_1_ready_to_source),
	.main_0_1_valid_from_source (auto_pthread_wrapper_inst_main_0_1_valid_from_source),
	.main_0_1_data_from_source (auto_pthread_wrapper_inst_main_0_1_data_from_source),
	.main_0_2_ready_from_sink (auto_pthread_wrapper_inst_main_0_2_ready_from_sink),
	.main_0_2_valid_to_sink (auto_pthread_wrapper_inst_main_0_2_valid_to_sink),
	.main_0_2_data_to_sink (auto_pthread_wrapper_inst_main_0_2_data_to_sink)
);



fwft_fifo main_0_2_inst (
	.clk (main_0_2_inst_clk),
	.reset (main_0_2_inst_reset),
	.clken (main_0_2_inst_clken),
	.write_en (main_0_2_inst_write_en),
	.write_data (main_0_2_inst_write_data),
	.read_en (main_0_2_inst_read_en),
	.read_data (main_0_2_inst_read_data),
	.full (main_0_2_inst_full),
	.almost_full (main_0_2_inst_almost_full),
	.empty (main_0_2_inst_empty),
	.almost_empty (main_0_2_inst_almost_empty),
	.usedw (main_0_2_inst_usedw)
);

defparam
	main_0_2_inst.width = 64,
	main_0_2_inst.depth = 10,
	main_0_2_inst.widthad = 4;


auto_pthread_wrapper_OC_1 auto_pthread_wrapper_OC_1_inst (
	.clk (auto_pthread_wrapper_OC_1_inst_clk),
	.reset (auto_pthread_wrapper_OC_1_inst_reset),
	.start (auto_pthread_wrapper_OC_1_inst_start),
	.finish (auto_pthread_wrapper_OC_1_inst_finish),
	.main_0_2_ready_to_source (auto_pthread_wrapper_OC_1_inst_main_0_2_ready_to_source),
	.main_0_2_valid_from_source (auto_pthread_wrapper_OC_1_inst_main_0_2_valid_from_source),
	.main_0_2_data_from_source (auto_pthread_wrapper_OC_1_inst_main_0_2_data_from_source),
	.main_0_3_ready_from_sink (auto_pthread_wrapper_OC_1_inst_main_0_3_ready_from_sink),
	.main_0_3_valid_to_sink (auto_pthread_wrapper_OC_1_inst_main_0_3_valid_to_sink),
	.main_0_3_data_to_sink (auto_pthread_wrapper_OC_1_inst_main_0_3_data_to_sink)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(*) begin
	main_inst_main_0_1_ready_from_sink = ~(main_0_1_inst_full);
end
always @(*) begin
	main_inst_main_0_3_valid_from_source = ~(main_0_3_inst_empty);
end
always @(*) begin
	main_inst_main_0_3_data_from_source = main_0_3_inst_read_data;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	main_0_1_inst_clk = clk;
end
always @(*) begin
	main_0_1_inst_reset = reset;
end
always @(*) begin
	main_0_1_inst_clken = ~(1'd0);
if (reset) begin main_0_1_inst_clken = 0; end
end
always @(*) begin
	main_0_1_inst_write_en = main_inst_main_0_1_valid_to_sink;
end
always @(*) begin
	main_0_1_inst_write_data = main_inst_main_0_1_data_to_sink;
end
always @(*) begin
	main_0_1_inst_read_en = auto_pthread_wrapper_inst_main_0_1_ready_to_source;
end
always @(*) begin
	main_0_3_inst_clk = clk;
end
always @(*) begin
	main_0_3_inst_reset = reset;
end
always @(*) begin
	main_0_3_inst_clken = ~(1'd0);
if (reset) begin main_0_3_inst_clken = 0; end
end
always @(*) begin
	main_0_3_inst_write_en = auto_pthread_wrapper_OC_1_inst_main_0_3_valid_to_sink;
end
always @(*) begin
	main_0_3_inst_write_data = auto_pthread_wrapper_OC_1_inst_main_0_3_data_to_sink;
end
always @(*) begin
	main_0_3_inst_read_en = main_inst_main_0_3_ready_to_source;
end
always @(*) begin
	auto_pthread_wrapper_inst_clk = clk;
end
always @(*) begin
	auto_pthread_wrapper_inst_reset = reset;
end
always @(*) begin
	auto_pthread_wrapper_inst_start = 1'd0;
	if ((main_inst_auto_pthread_wrapper_threadID == 16'd0)) begin
		auto_pthread_wrapper_inst_start = main_inst_auto_pthread_wrapper_start;
	end
end
always @(*) begin
	auto_pthread_wrapper_inst_main_0_1_valid_from_source = ~(main_0_1_inst_empty);
end
always @(*) begin
	auto_pthread_wrapper_inst_main_0_1_data_from_source = main_0_1_inst_read_data;
end
always @(*) begin
	auto_pthread_wrapper_inst_main_0_2_ready_from_sink = ~(main_0_2_inst_full);
end
always @(posedge clk) begin
	if ((reset | auto_pthread_wrapper_inst_start)) begin
		auto_pthread_wrapper_inst_finish_reg <= 1'd0;
	end
	if (auto_pthread_wrapper_inst_finish) begin
		auto_pthread_wrapper_inst_finish_reg <= 1'd1;
	end
end
always @(*) begin
	main_0_2_inst_clk = clk;
end
always @(*) begin
	main_0_2_inst_reset = reset;
end
always @(*) begin
	main_0_2_inst_clken = ~(1'd0);
if (reset) begin main_0_2_inst_clken = 0; end
end
always @(*) begin
	main_0_2_inst_write_en = auto_pthread_wrapper_inst_main_0_2_valid_to_sink;
end
always @(*) begin
	main_0_2_inst_write_data = auto_pthread_wrapper_inst_main_0_2_data_to_sink;
end
always @(*) begin
	main_0_2_inst_read_en = auto_pthread_wrapper_OC_1_inst_main_0_2_ready_to_source;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_clk = clk;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_reset = reset;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_start = 1'd0;
	if ((main_inst_auto_pthread_wrapper_OC_1_threadID == 16'd0)) begin
		auto_pthread_wrapper_OC_1_inst_start = main_inst_auto_pthread_wrapper_OC_1_start;
	end
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_main_0_2_valid_from_source = ~(main_0_2_inst_empty);
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_main_0_2_data_from_source = main_0_2_inst_read_data;
end
always @(*) begin
	auto_pthread_wrapper_OC_1_inst_main_0_3_ready_from_sink = ~(main_0_3_inst_full);
end
always @(posedge clk) begin
	if ((reset | auto_pthread_wrapper_OC_1_inst_start)) begin
		auto_pthread_wrapper_OC_1_inst_finish_reg <= 1'd0;
	end
	if (auto_pthread_wrapper_OC_1_inst_finish) begin
		auto_pthread_wrapper_OC_1_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	finish <= main_inst_finish;
end
always @(posedge clk) begin
	return_val <= main_inst_return_val;
end

endmodule
